`timescale 1ns/1ps
`include "config.vh"    // ADDR_WIDTH, PRI_BITS, K_LOG2, N_CORES

module gen_requests_k();
    // ---- Derived parameters ----
    localparam K_REQ = `K_LOG2;                    // requests per core
    localparam TOT_W = (1 + `ADDR_WIDTH + `PRI_BITS);

    // ---- Locals ----
    integer fd;
    integer c, i;
    integer seed;
    reg [`ADDR_WIDTH-1:0] addr;    // address field
    reg                   rw;      // 0=read, 1=write
    reg [`PRI_BITS-1:0]   prio;    // priority field
    reg [TOT_W-1:0]       packed;  // {rw, addr, prio}

    // File name as packed array (Vivado-friendly)
    reg [8*32-1:0] filename; // עד 32 תווים

    initial begin
        // Build file name for K_LOG2 up to 10
        if (`K_LOG2 < 10)
            filename = {"requests_K", "0"+`K_LOG2, ".mem"};
        else if (`K_LOG2 == 10)
            filename = {"requests_K10.mem"};
        else
            filename = {"requests_K", "X", ".mem"}; // fallback for unsupported

        // Open output file
        fd = $fopen(filename, "w");
        if (fd == 0) begin
            $display("ERROR: cannot open %0s for write.", filename);
            $finish;
        end

        // Header
        $fdisplay(fd, "// generated by gen_requests_k (pure Verilog)");
        $fdisplay(fd, "// K_LOG2=%0d, N_CORES=%0d, K_REQ=%0d, PRI_BITS=%0d, ADDR_WIDTH=%0d, TOT_W=%0d",
                      `K_LOG2, `N_CORES, K_REQ, `PRI_BITS, `ADDR_WIDTH, TOT_W);
        $fdisplay(fd, "// columns: core_index  request_index  packed_hex");

        // Generate requests
        seed = 32'h1234_5678;
        for (c = 0; c < `N_CORES; c = c + 1) begin
            seed = seed ^ (c * 32'h9E37_79B1);
            for (i = 0; i < K_REQ; i = i + 1) begin
                addr = $random(seed);
                rw   = $random(seed) & 1;
                prio = $random(seed) % (1 << `PRI_BITS);
                packed = {rw, addr, prio};
                $fdisplay(fd, "%0d %0d %0h", c, i, packed);
            end
        end

        $fclose(fd);
        $display("DONE: wrote %0d cores × %0d requests to %0s", `N_CORES, K_REQ, filename);
        $finish;
    end
endmodule
